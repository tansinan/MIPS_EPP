library ieee;
use ieee.std_logic_1164.all;

entity HighLatencyMathModule is
end entity;

architecture Behavioral of HighLatencyMathModule is
begin

end architecture;
