library ieee;
use ieee.std_logic_1164.all;

entity TypeRInstructionDecoder is
	instruction : in std_logic_vector(MIPS_CPU_INSTRUCTION_WIDTH - 1 downto 0);
end TypeRInstructionDecoder;

architecture Behavioral of TypeRInstructionDecoder is

begin


end Behavioral;

