library ieee;
use ieee.std_logic_1164.all;

entity TypeJInstructionDecoder is
	instruction : in std_logic_vector(MIPS_CPU_INSTRUCTION_WIDTH - 1 downto 0);
end TypeJInstructionDecoder;

architecture Behavioral of TypeJInstructionDecoder is

begin


end Behavioral;

