library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.MIPSCPU.all;

entity FlashRomController is
	port (
		clock: in Clock_t;
		reset: in Reset_t
	);
end entity;

architecture Behavioral of FlashRomController is
begin

end architecture;
