library ieee;
use ieee.std_logic_1164.all;

entity CP0PipelinePhaseInstructionDecode is
end entity;

architecture Behavioral of CP0PipelinePhaseInstructionDecode is
begin


end architecture;
