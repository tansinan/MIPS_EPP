library ieee;
use ieee.std_logic_1164.all;

entity CP0PipelinePhaseInstructionFetch is
end entity;

architecture Behavioral of CP0PipelinePhaseInstructionFetch is
begin


end architecture;

