library ieee;
use ieee.std_logic_1164.all;

package VirtualHardware is
	constant VIRTUAL_HARDWARE_RAM_FILE : string := "/mnt/MIPS_EPP_RAMDISK/RAM.txt";
	constant VIRTUAL_HARDWARE_RAM_TEMP_FILE : string := "/mnt/MIPS_EPP_RAMDISK/RAM_temp.txt";
end package;

package body VirtualHardware is
end package body;
