library ieee;
use ieee.std_logic_1164.all;
use work.MIPSCPU.all;
use work.MIPSCP0.all;

entity CP0Pipeline is
end entity;

architecture Behavioral of CP0Pipeline is
begin

end architecture;

