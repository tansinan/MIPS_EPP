library ieee;
use ieee.std_logic_1164.all;

entity PrimaryPipeline is
end entity;

architecture Behavioral of PrimaryPipeline is

begin


end architecture;

