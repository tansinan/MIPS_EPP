library ieee;
use ieee.std_logic_1164.all;

package MIPSCP0 is
	
end package;

package body MIPSCP0 is 
end package body;
