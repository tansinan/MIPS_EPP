library ieee;
use ieee.std_logic_1164.all;

entity CPOPipeline is
end CPOPipeline;

architecture Behavioral of CPOPipeline is
begin


end architecture;

