library ieee;
use ieee.std_logic_1164.all;

entity TypeIInstructionDecoder is
	instruction : in std_logic_vector(MIPS_CPU_INSTRUCTION_WIDTH - 1 downto 0);
end TypeIInstructionDecoder;

architecture Behavioral of TypeIInstructionDecoder is

begin


end Behavioral;

