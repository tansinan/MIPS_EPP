library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity PipelinePhaseExecute is
end PipelinePhaseExecute;

architecture Behavioral of PipelinePhaseExecute is

begin


end Behavioral;
