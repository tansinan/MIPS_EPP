library ieee;
use ieee.std_logic_1164.all;

entity HardwareRegisterMapper is
end entity;

architecture Behavioral of HardwareRegisterMapper is

begin


end architecture;

