library ieee;
use ieee.std_logic_1164.all;

entity CP0AddressTranslator is
end entity;

architecture Behavioral of CP0AddressTranslator is

begin


end architecture;

