library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity PipelinePhaseMemoryAccess is
end PipelinePhaseMemoryAccess;

architecture Behavioral of PipelinePhaseMemoryAccess is
begin


end Behavioral;
