library ieee;
use ieee.std_logic_1164.all;

entity PipelinePhaseWriteBack is
end PipelinePhaseWriteBack;

architecture Behavioral of PipelinePhaseWriteBack is

begin


end Behavioral;
